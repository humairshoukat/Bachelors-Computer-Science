module humairFADD(S,C,a,b,c);
input a,b,c;
output S,C;
wire axorb,ab,axorbc;
xor (axorb,a,b);
and (ab,a,b);
xor (S,axorb,c);
and (axorbc,axorb,c);
or (C,axorbc,ab);
endmodule

module test;
reg a,b,c;
wire S,C;
humairFADD x(S,C,a,b,c);
initial
begin
a=1'b 0; b=1'b 0; c=1'b 0;#10
a=1'b 0; b=1'b 0; c=1'b 1;#10
a=1'b 0; b=1'b 1; c=1'b 0;#10
a=1'b 0; b=1'b 1; c=1'b 1;#10
a=1'b 1; b=1'b 0; c=1'b 0;#10
a=1'b 1; b=1'b 0; c=1'b 1;#10
a=1'b 1; b=1'b 1; c=1'b 0;#10
a=1'b 1; b=1'b 1; c=1'b 1;#10
a=1'b 0; b=1'b 0; c=1'b 0;
end
endmodule
